//---------------------------------------------------------------------------------------------------//
// MIT License
//
// Copyright (c) 2022 José Luis Jiménez Arévalo, Eduardo García Olmos, Luis Alfredo Aceves Astengo
// 
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
// 
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
// 
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
//---------------------------------------------------------------------------------------------------//

module ram#(parameter DATA_SIZE=32,parameter SELEC_SIZE=16, parameter ADDRESSES=256)
	   (input logic clk,
	    input logic dm_we,
	    input logic [SELEC_SIZE-1:0] dm_address,
	    input logic [DATA_SIZE-1:0] dm_d,
	    output logic [DATA_SIZE-1:0] dm_q);
				
logic [DATA_SIZE-1:0] mem [ADDRESSES-1:0];
				
				
always_ff @(posedge clk) 
begin
	if (dm_we)
	begin
		mem[dm_address] <= dm_d;
	end
end
				
always_comb 
begin
	dm_q = mem[dm_address];
end

endmodule
